/home/tools/design_kits/cadence/GPDK045/gsclib045_svt_v4.4/gsclib045/lef/gsclib045_tech.lef